`timescale 1ns / 1ps


module mux_4x1_tb();
    reg [3:0] a;
    reg [1:0] s;
    wire o;
    
    mux_4x1 DUT(.i(a), .s(s), .F(o));
    
    initial begin
    
        s=0;
        a[0]=1 ; a[1]=0 ; a[2]=0 ; a[3]=0 ; #50 
        a[0]=0 ; a[1]=1 ; a[2]=0 ; a[3]=0 ; #50 
        a[0]=0 ; a[1]=0 ; a[2]=1 ; a[3]=0 ; #50 
        a[0]=0 ; a[1]=0 ; a[2]=0 ; a[3]=1 ; #50 
        
        s=1;
        a[0]=1 ; a[1]=0 ; a[2]=0 ; a[3]=0 ; #50 
        a[0]=0 ; a[1]=1 ; a[2]=0 ; a[3]=0 ; #50
        a[0]=0 ; a[1]=0 ; a[2]=1 ; a[3]=0 ; #50 
        a[0]=0 ; a[1]=0 ; a[2]=0 ; a[3]=1 ; #50 
        
        s=2;
        a[0]=1 ; a[1]=0 ; a[2]=0 ; a[3]=0 ; #50 
        a[0]=0 ; a[1]=1 ; a[2]=0 ; a[3]=0 ; #50 
        a[0]=0 ; a[1]=0 ; a[2]=1 ; a[3]=0 ; #50 
        a[0]=0 ; a[1]=0 ; a[2]=0 ; a[3]=1 ; #50 
        
        s=3;
        a[0]=1 ; a[1]=0 ; a[2]=0 ; a[3]=0 ; #50 
        a[0]=0 ; a[1]=1 ; a[2]=0 ; a[3]=0 ; #50 
        a[0]=0 ; a[1]=0 ; a[2]=1 ; a[3]=0 ; #50 
        a[0]=0 ; a[1]=0 ; a[2]=0 ; a[3]=1 ; #50 
        $finish();
    end
    
endmodule
